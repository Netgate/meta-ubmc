/*
 * Device Tree Source for AM33XX SoC
 *
 * Copyright (C) 2012 Texas Instruments Incorporated - http://www.ti.com/
 *
 * This file is licensed under the terms of the GNU General Public License
 * version 2.  This program is licensed "as is" without any warranty of any
 * kind, whether express or implied.
 */

#include <dt-bindings/gpio/gpio.h>
#include <dt-bindings/pinctrl/am33xx.h>

#include "skeleton.dtsi"

/ {
	compatible = "ti,am33xx";
	interrupt-parent = <&intc>;

	aliases {
		i2c0 = &i2c0;
		i2c1 = &i2c1;
		i2c2 = &i2c2;
		serial0 = &uart0;
		serial1 = &uart1;
		serial2 = &uart2;
		serial3 = &uart3;
		serial4 = &uart4;
		serial5 = &uart5;
		d_can0 = &dcan0;
		d_can1 = &dcan1;
		usb0 = &usb0;
		usb1 = &usb1;
		phy0 = &usb0_phy;
		phy1 = &usb1_phy;
		ethernet0 = &cpsw_emac0;
		ethernet1 = &cpsw_emac1;
	};

	cpus {
		#address-cells = <1>;
		#size-cells = <0>;
		cpu@0 {
			compatible = "arm,cortex-a8";
			device_type = "cpu";
			reg = <0>;

			/*
			 * To consider voltage drop between PMIC and SoC,
			 * tolerance value is reduced to 2% from 4% and
			 * voltage value is increased as a precaution.
			 */
			operating-points = <
				/* kHz    uV */
				720000  1285000
				600000  1225000
				500000  1125000
				275000  1125000
			>;
			voltage-tolerance = <2>; /* 2 percentage */

			clocks = <&dpll_mpu_ck>;
			clock-names = "cpu";

			clock-latency = <300000>; /* From omap-cpufreq driver */
		};
	};

	pmu {
		compatible = "arm,cortex-a8-pmu";
		interrupts = <3>;
	};

	/*
	 * The soc node represents the soc top level view. It is used for IPs
	 * that are not memory mapped in the MPU view or for the MPU itself.
	 */
	soc {
		compatible = "ti,omap-infra";
		mpu {
			compatible = "ti,omap3-mpu";
			ti,hwmods = "mpu";
		};
	};

	/*
	 * XXX: Use a flat representation of the AM33XX interconnect.
	 * The real AM33XX interconnect network is quite complex. Since
	 * it will not bring real advantage to represent that in DT
	 * for the moment, just use a fake OCP bus entry to represent
	 * the whole bus hierarchy.
	 */
	ocp {
		compatible = "simple-bus";
		#address-cells = <1>;
		#size-cells = <1>;
		ranges;
		ti,hwmods = "l3_main";

		l4_wkup: l4_wkup@44c00000 {
			compatible = "ti,am3-l4-wkup", "simple-bus";
			#address-cells = <1>;
			#size-cells = <1>;
			ranges = <0 0x44c00000 0x280000>;

			wkup_m3: wkup_m3@100000 {
				compatible = "ti,am3352-wkup-m3";
				reg = <0x100000 0x4000>,
				      <0x180000	0x2000>;
				reg-names = "umem", "dmem";
				ti,hwmods = "wkup_m3";
				ti,pm-firmware = "am335x-pm-firmware.elf";
			};

			prcm: prcm@200000 {
				compatible = "ti,am3-prcm";
				reg = <0x200000 0x4000>;

				prcm_clocks: clocks {
					#address-cells = <1>;
					#size-cells = <0>;
				};

				prcm_clockdomains: clockdomains {
				};
			};

			scm: scm@210000 {
				compatible = "ti,am3-scm", "simple-bus";
				reg = <0x210000 0x2000>;
				#address-cells = <1>;
				#size-cells = <1>;
				ranges = <0 0x210000 0x2000>;

				am33xx_pinmux: pinmux@800 {
					compatible = "pinctrl-single";
					reg = <0x800 0x238>;
					#address-cells = <1>;
					#size-cells = <0>;
					pinctrl-single,register-width = <32>;
					pinctrl-single,function-mask = <0x7f>;
				};

				scm_conf: scm_conf@0 {
					compatible = "syscon";
					reg = <0x0 0x800>;
					#address-cells = <1>;
					#size-cells = <1>;

					scm_clocks: clocks {
						#address-cells = <1>;
						#size-cells = <0>;
					};
				};

				wkup_m3_ipc: wkup_m3_ipc@1324 {
					compatible = "ti,am3352-wkup-m3-ipc";
					reg = <0x1324 0x24>;
					interrupts = <78>;
					ti,rproc = <&wkup_m3>;
					mboxes = <&mailbox &mbox_wkupm3>;
				};

				scm_clockdomains: clockdomains {
				};
			};
		};

		intc: interrupt-controller@48200000 {
			compatible = "ti,am33xx-intc";
			interrupt-controller;
			#interrupt-cells = <1>;
			reg = <0x48200000 0x1000>;
		};

		edma: edma@49000000 {
			compatible = "ti,edma3";
			ti,hwmods = "tpcc", "tptc0", "tptc1", "tptc2";
			reg =	<0x49000000 0x10000>,
				<0x44e10f90 0x40>;
			interrupts = <12 13 14>;
			#dma-cells = <1>;
		};

		gpio0: gpio@44e07000 {
			compatible = "ti,omap4-gpio";
			ti,hwmods = "gpio1";
			gpio-controller;
			#gpio-cells = <2>;
			interrupt-controller;
			#interrupt-cells = <2>;
			reg = <0x44e07000 0x1000>;
			interrupts = <96>;
		};

		gpio1: gpio@4804c000 {
			compatible = "ti,omap4-gpio";
			ti,hwmods = "gpio2";
			gpio-controller;
			#gpio-cells = <2>;
			interrupt-controller;
			#interrupt-cells = <2>;
			reg = <0x4804c000 0x1000>;
			interrupts = <98>;
		};

		gpio2: gpio@481ac000 {
			compatible = "ti,omap4-gpio";
			ti,hwmods = "gpio3";
			gpio-controller;
			#gpio-cells = <2>;
			interrupt-controller;
			#interrupt-cells = <2>;
			reg = <0x481ac000 0x1000>;
			interrupts = <32>;
		};

		gpio3: gpio@481ae000 {
			compatible = "ti,omap4-gpio";
			ti,hwmods = "gpio4";
			gpio-controller;
			#gpio-cells = <2>;
			interrupt-controller;
			#interrupt-cells = <2>;
			reg = <0x481ae000 0x1000>;
			interrupts = <62>;
		};

		uart0: serial@44e09000 {
			compatible = "ti,am3352-uart", "ti,omap3-uart";
			ti,hwmods = "uart1";
			clock-frequency = <48000000>;
			reg = <0x44e09000 0x2000>;
			interrupts = <72>;
			status = "disabled";
			dmas = <&edma 26>, <&edma 27>;
			dma-names = "tx", "rx";
		};

		uart1: serial@48022000 {
			compatible = "ti,am3352-uart", "ti,omap3-uart";
			ti,hwmods = "uart2";
			clock-frequency = <48000000>;
			reg = <0x48022000 0x2000>;
			interrupts = <73>;
			status = "disabled";
			dmas = <&edma 28>, <&edma 29>;
			dma-names = "tx", "rx";
		};

		uart2: serial@48024000 {
			compatible = "ti,am3352-uart", "ti,omap3-uart";
			ti,hwmods = "uart3";
			clock-frequency = <48000000>;
			reg = <0x48024000 0x2000>;
			interrupts = <74>;
			status = "disabled";
			dmas = <&edma 30>, <&edma 31>;
			dma-names = "tx", "rx";
		};

		uart3: serial@481a6000 {
			compatible = "ti,am3352-uart", "ti,omap3-uart";
			ti,hwmods = "uart4";
			clock-frequency = <48000000>;
			reg = <0x481a6000 0x2000>;
			interrupts = <44>;
			status = "disabled";
		};

		uart4: serial@481a8000 {
			compatible = "ti,am3352-uart", "ti,omap3-uart";
			ti,hwmods = "uart5";
			clock-frequency = <48000000>;
			reg = <0x481a8000 0x2000>;
			interrupts = <45>;
			status = "disabled";
		};

		uart5: serial@481aa000 {
			compatible = "ti,am3352-uart", "ti,omap3-uart";
			ti,hwmods = "uart6";
			clock-frequency = <48000000>;
			reg = <0x481aa000 0x2000>;
			interrupts = <46>;
			status = "disabled";
		};

		i2c0: i2c@44e0b000 {
			compatible = "ti,omap4-i2c";
			#address-cells = <1>;
			#size-cells = <0>;
			ti,hwmods = "i2c1";
			reg = <0x44e0b000 0x1000>;
			interrupts = <70>;
			status = "disabled";
		};

		i2c1: i2c@4802a000 {
			compatible = "ti,omap4-i2c";
			#address-cells = <1>;
			#size-cells = <0>;
			ti,hwmods = "i2c2";
			reg = <0x4802a000 0x1000>;
			interrupts = <71>;
			status = "disabled";
		};

		i2c2: i2c@4819c000 {
			compatible = "ti,omap4-i2c";
			#address-cells = <1>;
			#size-cells = <0>;
			ti,hwmods = "i2c3";
			reg = <0x4819c000 0x1000>;
			interrupts = <30>;
			status = "disabled";
		};

		mmc1: mmc@48060000 {
			compatible = "ti,omap4-hsmmc";
			ti,hwmods = "mmc1";
			ti,dual-volt;
			ti,needs-special-reset;
			ti,needs-special-hs-handling;
			dmas = <&edma 24
				&edma 25>;
			dma-names = "tx", "rx";
			interrupts = <64>;
			interrupt-parent = <&intc>;
			reg = <0x48060000 0x1000>;
			status = "disabled";
		};

		mmc2: mmc@481d8000 {
			compatible = "ti,omap4-hsmmc";
			ti,hwmods = "mmc2";
			ti,needs-special-reset;
			dmas = <&edma 2
				&edma 3>;
			dma-names = "tx", "rx";
			interrupts = <28>;
			interrupt-parent = <&intc>;
			reg = <0x481d8000 0x1000>;
			status = "disabled";
		};

		mmc3: mmc@47810000 {
			compatible = "ti,omap4-hsmmc";
			ti,hwmods = "mmc3";
			ti,needs-special-reset;
			interrupts = <29>;
			interrupt-parent = <&intc>;
			reg = <0x47810000 0x1000>;
			status = "disabled";
		};

		hwspinlock: spinlock@480ca000 {
			compatible = "ti,omap4-hwspinlock";
			reg = <0x480ca000 0x1000>;
			ti,hwmods = "spinlock";
			#hwlock-cells = <1>;
		};

		wdt2: wdt@44e35000 {
			compatible = "ti,omap3-wdt";
			ti,hwmods = "wd_timer2";
			reg = <0x44e35000 0x1000>;
			interrupts = <91>;
		};

		dcan0: can@481cc000 {
			compatible = "ti,am3352-d_can";
			ti,hwmods = "d_can0";
			reg = <0x481cc000 0x2000>;
			clocks = <&dcan0_fck>;
			clock-names = "fck";
			syscon-raminit = <&scm_conf 0x644 0>;
			interrupts = <52>;
			status = "disabled";
		};

		dcan1: can@481d0000 {
			compatible = "ti,am3352-d_can";
			ti,hwmods = "d_can1";
			reg = <0x481d0000 0x2000>;
			clocks = <&dcan1_fck>;
			clock-names = "fck";
			syscon-raminit = <&scm_conf 0x644 1>;
			interrupts = <55>;
			status = "disabled";
		};

		mailbox: mailbox@480C8000 {
			compatible = "ti,omap4-mailbox";
			reg = <0x480C8000 0x200>;
			interrupts = <77>;
			ti,hwmods = "mailbox";
			#mbox-cells = <1>;
			ti,mbox-num-users = <4>;
			ti,mbox-num-fifos = <8>;
			mbox_wkupm3: wkup_m3 {
				ti,mbox-tx = <0 0 0>;
				ti,mbox-rx = <0 0 3>;
			};
		};

		timer1: timer@44e31000 {
			compatible = "ti,am335x-timer-1ms";
			reg = <0x44e31000 0x400>;
			interrupts = <67>;
			ti,hwmods = "timer1";
			ti,timer-alwon;
		};

		timer2: timer@48040000 {
			compatible = "ti,am335x-timer";
			reg = <0x48040000 0x400>;
			interrupts = <68>;
			ti,hwmods = "timer2";
		};

		timer3: timer@48042000 {
			compatible = "ti,am335x-timer";
			reg = <0x48042000 0x400>;
			interrupts = <69>;
			ti,hwmods = "timer3";
		};

		timer4: timer@48044000 {
			compatible = "ti,am335x-timer";
			reg = <0x48044000 0x400>;
			interrupts = <92>;
			ti,hwmods = "timer4";
			ti,timer-pwm;
		};

		timer5: timer@48046000 {
			compatible = "ti,am335x-timer";
			reg = <0x48046000 0x400>;
			interrupts = <93>;
			ti,hwmods = "timer5";
			ti,timer-pwm;
		};

		timer6: timer@48048000 {
			compatible = "ti,am335x-timer";
			reg = <0x48048000 0x400>;
			interrupts = <94>;
			ti,hwmods = "timer6";
			ti,timer-pwm;
		};

		timer7: timer@4804a000 {
			compatible = "ti,am335x-timer";
			reg = <0x4804a000 0x400>;
			interrupts = <95>;
			ti,hwmods = "timer7";
			ti,timer-pwm;
		};

		usbotg_fck {
			#clock-cells = <0x0>;
			compatible = "ti,gate-clock";
			clocks = <0xb>;
			ti,bit-shift = <0x8>;
			reg = <0x47c>;
		};

		usb_tsc_fck {
			#clock-cells = <0x0>;
			compatible = "fixed-factor-clock";
			clocks = <0x5>;
			clock-mult = <0x1>;
			clock-div = <0x1>;
		};

		rtc: rtc@44e3e000 {
			compatible = "ti,am3352-rtc", "ti,da830-rtc";
			reg = <0x44e3e000 0x1000>;
			interrupts = <75
				      76>;
			ti,hwmods = "rtc";
		};

		spi0: spi@48030000 {
			compatible = "ti,omap4-mcspi";
			#address-cells = <1>;
			#size-cells = <0>;
			reg = <0x48030000 0x400>;
			interrupts = <65>;
			ti,spi-num-cs = <2>;
			ti,hwmods = "spi0";
			dmas = <&edma 16
				&edma 17
				&edma 18
				&edma 19>;
			dma-names = "tx0", "rx0", "tx1", "rx1";
			status = "disabled";
		};

		spi1: spi@481a0000 {
			compatible = "ti,omap4-mcspi";
			#address-cells = <1>;
			#size-cells = <0>;
			reg = <0x481a0000 0x400>;
			interrupts = <125>;
			ti,spi-num-cs = <2>;
			ti,hwmods = "spi1";
			dmas = <&edma 42
				&edma 43
				&edma 44
				&edma 45>;
			dma-names = "tx0", "rx0", "tx1", "rx1";
			status = "disabled";
		};

		usb: usb@47400000 {
			compatible = "ti,am33xx-usb";
			reg = <0x47400000 0x1000>;
			ranges;
			#address-cells = <1>;
			#size-cells = <1>;
			ti,hwmods = "usb_otg_hs";
			status = "okay";

			usb_ctrl_mod: control@44e10620 {
				compatible = "ti,am335x-usb-ctrl-module";
				reg = <0x44e10620 0x10
					0x44e10648 0x4>;
				reg-names = "phy_ctrl", "wakeup";
				status = "okay";
			};

			usb0_phy: usb-phy@47401300 {
				compatible = "ti,am335x-usb-phy";
				reg = <0x47401300 0x100>;
				reg-names = "phy";
				status = "okay";
				ti,ctrl_mod = <&usb_ctrl_mod>;
			};

			usb0: usb@47401000 {
				compatible = "ti,musb-am33xx";
				status = "okay";
				reg = <0x47401400 0x400
					0x47401000 0x200>;
				reg-names = "mc", "control";

				interrupts = <18>;
				interrupt-names = "mc";
				dr_mode = "host";
				mentor,multipoint = <1>;
				mentor,num-eps = <16>;
				mentor,ram-bits = <12>;
				mentor,power = <500>;
				phys = <&usb0_phy>;

				dmas = <&cppi41dma  0 0 &cppi41dma  1 0
					&cppi41dma  2 0 &cppi41dma  3 0
					&cppi41dma  4 0 &cppi41dma  5 0
					&cppi41dma  6 0 &cppi41dma  7 0
					&cppi41dma  8 0 &cppi41dma  9 0
					&cppi41dma 10 0 &cppi41dma 11 0
					&cppi41dma 12 0 &cppi41dma 13 0
					&cppi41dma 14 0 &cppi41dma  0 1
					&cppi41dma  1 1 &cppi41dma  2 1
					&cppi41dma  3 1 &cppi41dma  4 1
					&cppi41dma  5 1 &cppi41dma  6 1
					&cppi41dma  7 1 &cppi41dma  8 1
					&cppi41dma  9 1 &cppi41dma 10 1
					&cppi41dma 11 1 &cppi41dma 12 1
					&cppi41dma 13 1 &cppi41dma 14 1>;
				dma-names =
					"rx1", "rx2", "rx3", "rx4", "rx5", "rx6", "rx7",
					"rx8", "rx9", "rx10", "rx11", "rx12", "rx13",
					"rx14", "rx15",
					"tx1", "tx2", "tx3", "tx4", "tx5", "tx6", "tx7",
					"tx8", "tx9", "tx10", "tx11", "tx12", "tx13",
					"tx14", "tx15";
			};

			usb1_phy: usb-phy@47401b00 {
				compatible = "ti,am335x-usb-phy";
				reg = <0x47401b00 0x100>;
				reg-names = "phy";
				status = "okay";
				ti,ctrl_mod = <&usb_ctrl_mod>;
			};

			usb1: usb@47401800 {
				compatible = "ti,musb-am33xx";
				status = "okay";
				reg = <0x47401c00 0x400
					0x47401800 0x200>;
				reg-names = "mc", "control";
				interrupts = <19>;
				interrupt-names = "mc";
				dr_mode = "host";
				mentor,multipoint = <1>;
				mentor,num-eps = <10>;
				mentor,ram-bits = <12>;
				mentor,power = <500>;
				phys = <&usb1_phy>;

				dmas = <&cppi41dma 15 0 &cppi41dma 16 0
					&cppi41dma 17 0 &cppi41dma 18 0
					&cppi41dma 19 0 &cppi41dma 20 0
					&cppi41dma 21 0 &cppi41dma 22 0
					&cppi41dma 23 0 &cppi41dma 24 0
					&cppi41dma 25 0 &cppi41dma 26 0
					&cppi41dma 27 0 &cppi41dma 28 0
					&cppi41dma 29 0 &cppi41dma 15 1
					&cppi41dma 16 1 &cppi41dma 17 1
					&cppi41dma 18 1 &cppi41dma 19 1
					&cppi41dma 20 1 &cppi41dma 21 1
					&cppi41dma 22 1 &cppi41dma 23 1
					&cppi41dma 24 1 &cppi41dma 25 1
					&cppi41dma 26 1 &cppi41dma 27 1
					&cppi41dma 28 1 &cppi41dma 29 1>;
				dma-names =
					"rx1", "rx2", "rx3", "rx4", "rx5", "rx6", "rx7",
					"rx8", "rx9", "rx10", "rx11", "rx12", "rx13",
					"rx14", "rx15",
					"tx1", "tx2", "tx3", "tx4", "tx5", "tx6", "tx7",
					"tx8", "tx9", "tx10", "tx11", "tx12", "tx13",
					"tx14", "tx15";
			};

			cppi41dma: dma-controller@47402000 {
				compatible = "ti,am3359-cppi41";
				reg =  <0x47400000 0x1000
					0x47402000 0x1000
					0x47403000 0x1000
					0x47404000 0x4000>;
				reg-names = "glue", "controller", "scheduler", "queuemgr";
				interrupts = <17>;
				interrupt-names = "glue";
				#dma-cells = <2>;
				#dma-channels = <30>;
				#dma-requests = <256>;
				status = "disabled";
			};
		};

		epwmss0: epwmss@48300000 {
			compatible = "ti,am33xx-pwmss";
			reg = <0x48300000 0x10>;
			ti,hwmods = "epwmss0";
			#address-cells = <1>;
			#size-cells = <1>;
			status = "disabled";
			ranges = <0x48300100 0x48300100 0x80   /* ECAP */
				  0x48300180 0x48300180 0x80   /* EQEP */
				  0x48300200 0x48300200 0x80>; /* EHRPWM */

			ecap0: ecap@48300100 {
				compatible = "ti,am33xx-ecap";
				#pwm-cells = <3>;
				reg = <0x48300100 0x80>;
				interrupts = <31>;
				interrupt-names = "ecap0";
				ti,hwmods = "ecap0";
				status = "disabled";
			};

			ehrpwm0: ehrpwm@48300200 {
				compatible = "ti,am33xx-ehrpwm";
				#pwm-cells = <3>;
				reg = <0x48300200 0x80>;
				ti,hwmods = "ehrpwm0";
				status = "disabled";
			};
		};

		epwmss1: epwmss@48302000 {
			compatible = "ti,am33xx-pwmss";
			reg = <0x48302000 0x10>;
			ti,hwmods = "epwmss1";
			#address-cells = <1>;
			#size-cells = <1>;
			status = "disabled";
			ranges = <0x48302100 0x48302100 0x80   /* ECAP */
				  0x48302180 0x48302180 0x80   /* EQEP */
				  0x48302200 0x48302200 0x80>; /* EHRPWM */

			ecap1: ecap@48302100 {
				compatible = "ti,am33xx-ecap";
				#pwm-cells = <3>;
				reg = <0x48302100 0x80>;
				interrupts = <47>;
				interrupt-names = "ecap1";
				ti,hwmods = "ecap1";
				status = "disabled";
			};

			ehrpwm1: ehrpwm@48302200 {
				compatible = "ti,am33xx-ehrpwm";
				#pwm-cells = <3>;
				reg = <0x48302200 0x80>;
				ti,hwmods = "ehrpwm1";
				status = "disabled";
			};
		};

		epwmss2: epwmss@48304000 {
			compatible = "ti,am33xx-pwmss";
			reg = <0x48304000 0x10>;
			ti,hwmods = "epwmss2";
			#address-cells = <1>;
			#size-cells = <1>;
			status = "disabled";
			ranges = <0x48304100 0x48304100 0x80   /* ECAP */
				  0x48304180 0x48304180 0x80   /* EQEP */
				  0x48304200 0x48304200 0x80>; /* EHRPWM */

			ecap2: ecap@48304100 {
				compatible = "ti,am33xx-ecap";
				#pwm-cells = <3>;
				reg = <0x48304100 0x80>;
				interrupts = <61>;
				interrupt-names = "ecap2";
				ti,hwmods = "ecap2";
				status = "disabled";
			};

			ehrpwm2: ehrpwm@48304200 {
				compatible = "ti,am33xx-ehrpwm";
				#pwm-cells = <3>;
				reg = <0x48304200 0x80>;
				ti,hwmods = "ehrpwm2";
				status = "disabled";
			};
		};

		mac: ethernet@4a100000 {
			compatible = "ti,am335x-cpsw","ti,cpsw";
			ti,hwmods = "cpgmac0";
			clocks = <&cpsw_125mhz_gclk>, <&cpsw_cpts_rft_clk>;
			clock-names = "fck", "cpts";
			cpdma_channels = <8>;
			ale_entries = <1024>;
			bd_ram_size = <0x2000>;
			no_bd_ram = <0>;
			rx_descs = <64>;
			mac_control = <0x20>;
			slaves = <2>;
			active_slave = <0>;
			cpts_clock_mult = <0x80000000>;
			cpts_clock_shift = <29>;
			reg = <0x4a100000 0x800
			       0x4a101200 0x100>;
			#address-cells = <1>;
			#size-cells = <1>;
			interrupt-parent = <&intc>;
			/*
			 * c0_rx_thresh_pend
			 * c0_rx_pend
			 * c0_tx_pend
			 * c0_misc_pend
			 */
			interrupts = <40 41 42 43>;
			ranges;
			syscon = <&scm_conf>;
			status = "disabled";

			davinci_mdio: mdio@4a101000 {
				compatible = "ti,davinci_mdio";
				#address-cells = <1>;
				#size-cells = <0>;
				ti,hwmods = "davinci_mdio";
				bus_freq = <1000000>;
				reg = <0x4a101000 0x100>;
				status = "disabled";
			};

			cpsw_emac0: slave@4a100200 {
				/* Filled in by U-Boot */
				mac-address = [ 00 00 00 00 00 00 ];
			};

			cpsw_emac1: slave@4a100300 {
				/* Filled in by U-Boot */
				mac-address = [ 00 00 00 00 00 00 ];
			};

			phy_sel: cpsw-phy-sel@44e10650 {
				compatible = "ti,am3352-cpsw-phy-sel";
				reg= <0x44e10650 0x4>;
				reg-names = "gmii-sel";
			};
		};

		ocmcram: ocmcram@40300000 {
			compatible = "mmio-sram";
			reg = <0x40300000 0x10000>; /* 64k */
		};

		elm: elm@48080000 {
			compatible = "ti,am3352-elm";
			reg = <0x48080000 0x2000>;
			interrupts = <4>;
			ti,hwmods = "elm";
			status = "disabled";
		};

		lcdc: lcdc@4830e000 {
			compatible = "ti,am33xx-tilcdc";
			reg = <0x4830e000 0x1000>;
			interrupt-parent = <&intc>;
			interrupts = <36>;
			ti,hwmods = "lcdc";
			status = "disabled";
		};

		tscadc: tscadc@44e0d000 {
			compatible = "ti,am3359-tscadc";
			reg = <0x44e0d000 0x1000>;
			interrupt-parent = <0x1>;
			interrupts = <0x10>;
			ti,hwmods = "adc_tsc";
			status = "okay";

			tsc {
				compatible = "ti,am3359-tsc";
				ti,wires = <0x4>;
				ti,x-plate-resistance = <0xc8>;
				ti,coordinate-readouts = <0x5>;
				ti,wire-config = <0x0 0x11 0x22 0x33>;
				ti,charge-delay = <0x400>;
			};

			adc {
				#io-channel-cells = <0x1>;
				compatible = "ti,am3359-adc";
				ti,adc-channels = <0x4 0x5 0x6 0x7>;
			};
		};

		gpmc: gpmc@50000000 {
			compatible = "ti,am3352-gpmc";
			ti,hwmods = "gpmc";
			ti,no-idle-on-init;
			reg = <0x50000000 0x2000>;
			interrupts = <100>;
			gpmc,num-cs = <7>;
			gpmc,num-waitpins = <2>;
			#address-cells = <2>;
			#size-cells = <1>;
			status = "disabled";
		};

		sham: sham@53100000 {
			compatible = "ti,omap4-sham";
			ti,hwmods = "sham";
			reg = <0x53100000 0x200>;
			interrupts = <109>;
			dmas = <&edma 36>;
			dma-names = "rx";
		};

		aes: aes@53500000 {
			compatible = "ti,omap4-aes";
			ti,hwmods = "aes";
			reg = <0x53500000 0xa0>;
			interrupts = <103>;
			dmas = <&edma 6>,
			       <&edma 5>;
			dma-names = "tx", "rx";
		};

		mcasp0: mcasp@48038000 {
			compatible = "ti,am33xx-mcasp-audio";
			ti,hwmods = "mcasp0";
			reg = <0x48038000 0x2000>,
			      <0x46000000 0x400000>;
			reg-names = "mpu", "dat";
			interrupts = <80>, <81>;
			interrupt-names = "tx", "rx";
			status = "disabled";
			dmas = <&edma 8>,
				<&edma 9>;
			dma-names = "tx", "rx";
		};

		mcasp1: mcasp@4803C000 {
			compatible = "ti,am33xx-mcasp-audio";
			ti,hwmods = "mcasp1";
			reg = <0x4803C000 0x2000>,
			      <0x46400000 0x400000>;
			reg-names = "mpu", "dat";
			interrupts = <82>, <83>;
			interrupt-names = "tx", "rx";
			status = "disabled";
			dmas = <&edma 10>,
				<&edma 11>;
			dma-names = "tx", "rx";
		};

		rng: rng@48310000 {
			compatible = "ti,omap4-rng";
			ti,hwmods = "rng";
			reg = <0x48310000 0x2000>;
			interrupts = <111>;
		};
	};
};

/include/ "am33xx-clocks.dtsi"
